`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 02/20/2020 12:07:34 PM
// Design Name: 
// Module Name: charROM
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module charROM(
    input [6:0] addr,
    output reg [63:0] data 
);
    
    always @(*) begin
        case(addr)
            7'd0:   data = 64'h0000000000000000;
            7'd1:   data = 64'h0000000000000000;
            7'd2:   data = 64'h0000000000000000;
            7'd3:   data = 64'h0000000000000000;
            7'd4:   data = 64'h0000000000000000;
            7'd5:   data = 64'h0000000000000000;
            7'd6:   data = 64'h0000000000000000;
            7'd7:   data = 64'h0000000000000000;
            7'd8:   data = 64'h0000000000000000;
            7'd9:   data = 64'h0000000000000000;
            7'd10:  data = 64'h0000000000000000;
            7'd11:  data = 64'h0000000000000000;
            7'd12:  data = 64'h0000000000000000;
            7'd13:  data = 64'h0000000000000000;
            7'd14:  data = 64'h0000000000000000;
            7'd15:  data = 64'h0000000000000000;
            7'd16:  data = 64'h0000000000000000;
            7'd17:  data = 64'h0000000000000000;
            7'd18:  data = 64'h0000000000000000;
            7'd19:  data = 64'h0000000000000000;
            7'd20:  data = 64'h0000000000000000;
            7'd21:  data = 64'h0000000000000000;
            7'd22:  data = 64'h0000000000000000;
            7'd23:  data = 64'h0000000000000000;
            7'd24:  data = 64'h0000000000000000;
            7'd25:  data = 64'h0000000000000000;
            7'd26:  data = 64'h0000000000000000;
            7'd27:  data = 64'h0000000000000000;
            7'd28:  data = 64'h0000000000000000;
            7'd29:  data = 64'h0000000000000000;
            7'd30:  data = 64'h0000000000000000;
            7'd31:  data = 64'h0000000000000000;
            7'd32:  data = 64'h0000000000000000;
            7'd33:  data = 64'h0000005f00000000;
            7'd34:  data = 64'h0000030003000000;
            7'd35:  data = 64'h643c26643c262400;
            7'd36:  data = 64'h2649497f49493200;
            7'd37:  data = 64'h4225120824522100;
            7'd38:  data = 64'h20504e5522582800;
            7'd39:  data = 64'h0000000300000000;
            7'd40:  data = 64'h00001c2241000000;
            7'd41:  data = 64'h00000041221c0000;
            7'd42:  data = 64'h0015150e0e151500;
            7'd43:  data = 64'h0008083e08080000;
            7'd44:  data = 64'h0000005030000000;
            7'd45:  data = 64'h0008080808080000;
            7'd46:  data = 64'h0000004000000000;
            7'd47:  data = 64'h4020100804020100;
            7'd48:  data = 64'h003e4141413e0000;
            7'd49:  data = 64'h0000417f40000000;
            7'd50:  data = 64'h00426151496e0000;
            7'd51:  data = 64'h0022414949360000;
            7'd52:  data = 64'h001814127f100000;
            7'd53:  data = 64'h0027494949710000;
            7'd54:  data = 64'h003c4a4948700000;
            7'd55:  data = 64'h004321110d030000;
            7'd56:  data = 64'h0036494949360000;
            7'd57:  data = 64'h00060949291e0000;
            7'd58:  data = 64'h0000001200000000;
            7'd59:  data = 64'h0000005230000000;
            7'd60:  data = 64'h0000081414220000;
            7'd61:  data = 64'h0014141414141400;
            7'd62:  data = 64'h0000221414080000;
            7'd63:  data = 64'h0002015905020000;
            7'd64:  data = 64'h3e415d554d512e00;
            7'd65:  data = 64'h407c4a094a7c4000; //A
            7'd66:  data = 64'h417f494949493600; //B
            7'd67:  data = 64'h1c22414141412200; //C
            7'd68:  data = 64'h417f414141221c00;
            7'd69:  data = 64'h417f49495d416300;
            7'd70:  data = 64'h417f49091d010300;
            7'd71:  data = 64'h1c224149493a0800;
            7'd72:  data = 64'h417f0808087f4100;
            7'd73:  data = 64'h0041417F41410000;
            7'd74:  data = 64'h304041413F010100;
            7'd75:  data = 64'h417f080c12614100;
            7'd76:  data = 64'h417f414040406000;
            7'd77:  data = 64'h417f420c427f4100;
            7'd78:  data = 64'h417f420c117f0100;
            7'd79:  data = 64'h1c22414141221c00;
            7'd80:  data = 64'h417f490909090600;
            7'd81:  data = 64'h0c12212161524c00;
            7'd82:  data = 64'h417f090919694600;
            7'd83:  data = 64'h6649494949493300;
            7'd84:  data = 64'h0301417f41010300;
            7'd85:  data = 64'h013f4140413f0100;
            7'd86:  data = 64'h010f3140310f0100;
            7'd87:  data = 64'h011f6114611f0100;
            7'd88:  data = 64'h4141360836414100;
            7'd89:  data = 64'h0103447844030100;
            7'd90:  data = 64'h4361514945436100;
            7'd91:  data = 64'h00007f4141000000;
            7'd92:  data = 64'h0102040810204000;
            7'd93:  data = 64'h000041417f000000;
            7'd94:  data = 64'h0004020101020400;
            7'd95:  data = 64'h0040404040404000;
            7'd96:  data = 64'h0001020000000000;
            7'd97:  data = 64'h00344a4a4a3c4000;
            7'd98:  data = 64'h00413f4848483000;
            7'd99:  data = 64'h003c424242240000;
            7'd100: data = 64'h00304848493f4000;
            7'd101: data = 64'h003c4a4a4a2c0000;
            7'd102: data = 64'h0000487e49090000;
            7'd103: data = 64'h00264949493f0100;
            7'd104: data = 64'h417f480444784000;
            7'd105: data = 64'h0000447d40000000;
            7'd106: data = 64'h000040443d000000;
            7'd107: data = 64'h417f101824424200;
            7'd108: data = 64'h0040417f40400000;
            7'd109: data = 64'h427e027c027e4000;
            7'd110: data = 64'h427e4402427c4000;
            7'd111: data = 64'h003c4242423c0000;
            7'd112: data = 64'h00417f4909090600;
            7'd113: data = 64'h00060909497f4100;
            7'd114: data = 64'h00427e4402020400;
            7'd115: data = 64'h00644a4a4a360000;
            7'd116: data = 64'h00043f4444200000;
            7'd117: data = 64'h00023e4040227e40;
            7'd118: data = 64'h020e3240320e0200;
            7'd119: data = 64'h021e6218621e0200;
            7'd120: data = 64'h4262140814624200;
            7'd121: data = 64'h0143453805030100;
            7'd122: data = 64'h004662524a466200;
            7'd123: data = 64'h0000083641000000;
            7'd124: data = 64'h0000007f00000000;
            7'd125: data = 64'h0000004136080000;
            7'd126: data = 64'h0018080810101800;
            7'd127: data = 64'hAA55AA55AA55AA55;
            default: data = 64'h0000000000000000;
        endcase
    end
    
endmodule